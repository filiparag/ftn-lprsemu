------------------------------------------------------------------
        "000000000000000";
end architecture;
