------------------------------------------------------------------

	oQ <= rMEM(to_integer(unsigned(iA)));

end architecture;
